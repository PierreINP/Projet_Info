--commentaire
library ieee; --use lib
--a virer s<= a+b;
